// AHBGPIO testbench

program automatic AHBGPIO_tb
    (AHBGPIO_intf.DRIVER ahbgpio_intf);


// Test bench
    initial 
    begin 


    end

endprogram