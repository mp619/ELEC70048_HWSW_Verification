module multiplier_stim ();


    
endmodule